11110110101010111010001101100110110011011000001010110111100100001111010110011100111101100001011001101100000100101_0000000000000000000000000000000000000000000000000000000000000000000000000000																							
01110100011010001011011000000100011011011000101010101000000000100101100001100101011100110011001111110111011010100_1101010101110100011011001101100110110000010111101100001011001101100000100101																							
00111011001000101010010100010000100100001100101011111111000011001000011000101111101101000011111111100111001100100_1101110101110100011011001101100110110000010101101111001000011110101100111001																							
11110100001000011001100001111110010101010111111010111010111100001110000001011011011000001110110110101101001001100_0100110100010110110000001000110110110001010111100110011001111110111011010100																							
00111000000001000000110001100101011111101000001010101011110011111010001101010011111111001011110110100001000000101_1101010100010110110000001000110110110001010101010000000001001011000011001010																							
00110110100010000011000101011000001111010111101010000000001010100000100110101111010000010101100110100100101010010_0110010001010100101000100001001000011001010101101000011111111100111001100100																							
01110000100101001000101011001010110001101001000011110100110110101100110001110111000100100101000010101100100100010_0110110001010100101000100001001000011001010111111110000110010000110001011111																							
11111000101010001010001100000011001101000101110011000001001011111000100010011101111100011011101011011010001110101_1100010000110011000011111100101010101111110111000001110110110101101001001100																							
10110000101101111010100010011100101110000010000010101010110111100100001100101000000010101000010110001011011000110_1101010000110011000011111100101010101111110101110101111000011100000010110110																							
00111011011011100111001010100010001111000110100010001001110000111111010001011110010111011010110000101101110000011_0100000010000001100011001010111111010000010111111001011110110100001000000101																							