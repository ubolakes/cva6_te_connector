11110110101010110100011001101001101000000111110011010000100100110010110101010010110001110111100001011011110110101_0000000000000000000000000000000000000000000000000000000000000000000000000000																							
01110100011010000010110001101100111011100001111010100001011010101000100000011110110010100110001010101000111100110_1101010101101000110011010011010000001111100110001110111100001011011110110101																							
00111011001000111011011010011000111011001100111010011011001011100100100001000111011110111110111010001111001010000_1101110101101000110011010011010000001111100110100001001001100101101010100101																							
11110100001000010011000110101101001001010111010011001111101000111010100101011000100100100110100001001000011111101_1100110100000101100011011001110111000011110110010100110001010101000111100110																							
00111000000001000101001100101001000011111110111010001010010100110100101000001011000000110001000101011010111011100_0101010100000101100011011001110111000011110101000010110101010001000000111101																							
00110110100010010101110111111101000010011010100010001100110111101001001111111101111100101111011110111011101001010_1100010000100110001101011010010010101110100100100100110100001001000011111101																							
01110000100101000101000100111000101010010011101010011010101011111101111010010000101101010100111010111100110111101_1101010000100110001101011010010010101110100110011111010001110101001010110001																							
11111000101010000100011011110110101110000001100010010110110010100011011010110000101000010100001110000010111110000_1101001010001010001001110001010100100111010101101010100111010111100110111101																							
10110000101101110001000010000111111110000010111011000100010110000010000011000010011111111101001000011001001111011_0100001010001010001001110001010100100111010100110101010111111011110100100001																							
00111011011011100101000110111100111101100000110011001010111011101000000010111101011001000000000101101000001101101_1101010100001000110111101101011100000011000101000010100001110000010111110000