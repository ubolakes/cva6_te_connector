11110110101010101001101000111011001110010100110010111100011100100111000100010001111000000000000100000010001101101_1101110101010011010001110110011100101001100101111000111001001110001000100011
01110100011010010000010001010011010010010000111010000101010101110101110110000100011100011111000001111110001010111_1101010100010011010001110110011100101001100111000000000000100000010001101101
00111011001000110011010110101011111000111000011011101100010110000100010000110100111010100100011110010010010010000_0101010001100000100010100110100100100001110100001010101011101011101100001000
11110100001000010011011101100101100010010010011011001110101101000110110101111010110001111010110011010011011110010_1100110000100000100010100110100100100001110111100011111000001111110001010111
00111000000001000110000011010010011000010001010010011101110010011111111111111110111000111010001101101111000100100_0110100010100110101101010111110001110000110111011000101100001000100001101001
00110110100010011101100000110101110010100001111010100010010001010111010001000100110001100010101001001110001100001_0110000100100110101101010111110001110000110111010100100011110010010010010000
01110000100101011001000110110001000000100101000010100110011011111001011110110000001001101100100000100001010111101_1101001010100110111011001011000100100100110110011101011010001101101011110101
11111000101010000110101010110110010101100100111011110001111010100011100011110011011000110011100011010100110100110_1100010100100110111011001011000100100100110110001111010110011010011011110010
10110000101101100010010100001110101101010001111011010101100001100000111100110001001001101111001011100111111001101_0110011011001100000110100100110000100010100100111011100100111111111111111101